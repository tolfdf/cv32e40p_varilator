module test_pkg_import;
  import perturbation_pkg::*;
endmodule
